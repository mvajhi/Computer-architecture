module data_path(
    input pcsel,
    input regsel,
    input extend_func,
    input wereg,
    input wedata,
    input aluselb,
    input aluop,
    input outsel,
    output op,
    output func3,
    output func7
);

endmodule