module adder(
    input [31:0] A,
    input [31:0] B,
    output [31:0] C,
    output reg co
);
    assign {co, C} = A + B;
endmodule
